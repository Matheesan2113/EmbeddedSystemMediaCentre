-- Implements a simple Nios II system for the DE2 board.
-- Inputs: SW7-0 are parallel port inputs to the Nios II system.
-- CLOCK_50 is the system clock.
-- KEY0 is the active-low system reset.
-- Outputs: LEDG7-0 are parallel port outputs from the Nios II system.
-- SDRAM ports correspond to the signals in Figure 2; their names are those
-- used in the DE2 User Manual.
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY System2 IS
	PORT ( 
		SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		CLOCK_50 : IN STD_LOGIC;
		LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		LCD_EN : OUT STD_LOGIC;
		LCD_RW : OUT STD_LOGIC;
		LCD_RS : OUT STD_LOGIC;
		LCD_ON : OUT STD_LOGIC;
		LCD_DATA: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
		DRAM_ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		DRAM_BA_1, DRAM_BA_0 : BUFFER STD_LOGIC;
		DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
		DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		DRAM_UDQM, DRAM_LDQM : BUFFER STD_LOGIC );
		
END System2;

ARCHITECTURE Structure OF System2 IS

COMPONENT nios_system
	PORT ( 
		clk : IN STD_LOGIC;
		reset_n : IN STD_LOGIC;
		out_port_from_the_LEDs : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		in_port_to_the_Switches : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		
		-- the_lcd_16207_0
        LCD_E_from_the_lcd_16207_0 : OUT STD_LOGIC;
        LCD_RS_from_the_lcd_16207_0 : OUT STD_LOGIC;
        LCD_RW_from_the_lcd_16207_0 : OUT STD_LOGIC;
        LCD_data_to_and_from_the_lcd_16207_0 : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

		zs_addr_from_the_sdram: OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		zs_ba_from_the_sdram: BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
		zs_cas_n_from_the_sdram: OUT STD_LOGIC;
		zs_cke_from_the_sdram: OUT STD_LOGIC;
		zs_cs_n_from_the_sdram: OUT STD_LOGIC;
		zs_dq_to_and_from_the_sdram: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		zs_dqm_from_the_sdram: BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
		zs_ras_n_from_the_sdram: OUT STD_LOGIC;
		zs_we_n_from_the_sdram: OUT STD_LOGIC );
END COMPONENT;

COMPONENT sdram_pll
	PORT ( 
		inclk0 : IN STD_LOGIC;
		c0 : OUT STD_LOGIC );
END COMPONENT;

SIGNAL BA : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL DQM : STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN
	--BA <= (DRAM_BA_1 & DRAM_BA_0);
	--DQM <= (DRAM_UDQM & DRAM_LDQM);
	DRAM_BA_1 <= BA(1);
	DRAM_BA_0 <= BA(0);
	
	DRAM_UDQM <= DQM(1);
	DRAM_LDQM <= DQM(0);
	
	-- Instantiate the Nios II system entity generated by the SOPC Builder.
	NiosII: nios_system PORT MAP (CLOCK_50, '1', LEDG, SW, LCD_EN, LCD_RS, LCD_RW, LCD_DATA,
								DRAM_ADDR, BA, DRAM_CAS_N, DRAM_CKE, DRAM_CS_N,
								DRAM_DQ, DQM, DRAM_RAS_N, DRAM_WE_N );
	
	-- Instantiate the entity sdram_pll (inclk0, c0).
	neg_3ns: sdram_pll PORT MAP (CLOCK_50, DRAM_CLK);
	LCD_ON <= '1';
END Structure;